
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity seven_segment_timer is
Port ( );
end seven_segment_timer;

architecture Behavioral of seven_segment_timer is

begin


end Behavioral;
